LIBRARY ieee;
USE ieee.std_logic_1164.all;


ENTITY airplane_cl is
	PORT(clock, resetn, ivalid, iready: IN std_logic;
		  datain: IN std_logic_vector(7 downto 0);
		  oready, ovalid: OUT std_logic;
		  dataout: OUT std_logic_vector(7 downto 0));
END airplane_cl;

ARCHITECTURE structure of airplane_cl is
	--Declare the component, then port map it!

	BEGIN


END structure;
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
	
	
	

/////////////////////////////////////////////////////////////////
// MODULE mat_cl_system
/////////////////////////////////////////////////////////////////
module mat_cl_system
(
   input logic clock,
   input logic clock2x,
   input logic resetn
);
endmodule

